----------------------------------------------------------------------------------
-- utils_pkg.vhdl
--
-- Description: defines some common macros and functions
----------------------------------------------------------------------------------

-- utils_pkg.vhdl

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

----------------------------------------------------------------------------------
-- Package header
----------------------------------------------------------------------------------

package utils_pkg is

    constant DATA_WIDTH : integer := 32;

end package utils_pkg;
